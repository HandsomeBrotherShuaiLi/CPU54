`timescale 1ns / 1ps

module Reg_DMUX(
    input [4:0] iData,
    input iEna,
    output reg [31:0] oData
    );
    always @(*)
    begin
    if(iEna==1)
    begin
    case(iData)
    5'b00000:oData=32'b00000000_00000000_00000000_00000001;
    5'b00001:oData=32'b00000000_00000000_00000000_00000010;
    5'b00010:oData=32'b00000000_00000000_00000000_00000100;
    5'b00011:oData=32'b00000000_00000000_00000000_00001000;
    5'b00100:oData=32'b00000000_00000000_00000000_00010000;
    5'b00101:oData=32'b00000000_00000000_00000000_00100000;
    5'b00110:oData=32'b00000000_00000000_00000000_01000000;
    5'b00111:oData=32'b00000000_00000000_00000000_10000000;
    //8
    5'b01000:oData=32'b00000000_00000000_00000001_00000000;
    5'b01001:oData=32'b00000000_00000000_00000010_00000000;
    5'b01010:oData=32'b00000000_00000000_00000100_00000000;
    5'b01011:oData=32'b00000000_00000000_00001000_00000000;
    5'b01100:oData=32'b00000000_00000000_00010000_00000000;
    5'b01101:oData=32'b00000000_00000000_00100000_00000000;
    5'b01110:oData=32'b00000000_00000000_01000000_00000000;
    5'b01111:oData=32'b00000000_00000000_10000000_00000000;
    //16
    5'b10000:oData=32'b00000000_00000001_00000000_00000000;
    5'b10001:oData=32'b00000000_00000010_00000000_00000000;
    5'b10010:oData=32'b00000000_00000100_00000000_00000000;
    5'b10011:oData=32'b00000000_00001000_00000000_00000000;
    5'b10100:oData=32'b00000000_00010000_00000000_00000000;
    5'b10101:oData=32'b00000000_00100000_00000000_00000000;
    5'b10110:oData=32'b00000000_01000000_00000000_00000000;
    5'b10111:oData=32'b00000000_10000000_00000000_00000000;
    //24
    5'b11000:oData=32'b00000001_00000000_00000000_00000000;
    5'b11001:oData=32'b00000010_00000000_00000000_00000000;
    5'b11010:oData=32'b00000100_00000000_00000000_00000000;
    5'b11011:oData=32'b00001000_00000000_00000000_00000000;
    5'b11100:oData=32'b00010000_00000000_00000000_00000000;
    5'b11101:oData=32'b00100000_00000000_00000000_00000000;
    5'b11110:oData=32'b01000000_00000000_00000000_00000000;
    5'b11111:oData=32'b10000000_00000000_00000000_00000000;
    //32
    endcase
    end
    else
      begin
      oData=32'b00000000_00000000_00000000_00000000;
      end
    end
endmodule